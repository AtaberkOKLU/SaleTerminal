
module FP_MULT (
	dataa,
	datab,
	n,
	result);	

	input	[31:0]	dataa;
	input	[31:0]	datab;
	input	[3:0]	n;
	output	[31:0]	result;
endmodule
